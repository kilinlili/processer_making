module mem1(
    output [1:0] fromP_SIZE,
    output fromP_MEMWRITE,fromP_MEMREAD,
    output [31:0] toADDRESS,WRITEDATA,
    input[31:0] LOADDATA
);

endmodule 